library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity top is

port (

);

end;
architecture behaviour of top is

begin


end architecture;
